module Digital_Clock;


endmodule