module UART_Transmitter
(
    output wire dout,
    input wire [7:0] data,
    input wire start,
    input wire dnum,snum,
    input wire [1:0] bd_rate,par,
    input wire clk,rst,en
);


// declaring signals




// binary counter






endmodule