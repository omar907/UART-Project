module Baudrate_Generator;


endmodule