 module UART_Receiver
 (
    input wire data_bit,
    output wire [7:0] data
 );
 
 
 endmodule