 module UART_Receiver
 (
    input wire din,
    input wire dnum,snum,
    input wire bd_rate,par,
    
    input clk,rst,
    
    output wire [7:0] data,
    output error
 );
 
 
 
 
 
 endmodule